module HiCore_cmt_branch(
    
)